--FUNDUMENTAL CELL - METHODE I:
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RCPFA_CELL_I IS
    PORT(
        A, B : IN STD_LOGIC;
        FIN, CIN : IN STD_LOGIC;
        FOUT, COUT: OUT STD_LOGIC;
        S : OUT STD_LOGIC
    );
END ENTITY RCPFA_CELL_I;
ARCHITECTURE RCPFA_CELL_I_ARC OF RCPFA_CELL_I IS
    SIGNAL Y : STD_LOGIC;
BEGIN
    FOUT <= NOT (A NAND B);
    Y <= (A OR B) NAND (NOT CIN);
    S <= Y NAND (NOT FIN);
    COUT <= NOT(Y NAND NOT(NOT FIN));
END ARCHITECTURE RCPFA_CELL_I_ARC;
-----------------------------------------------------------------------------------
--FUNDUMENTAL CELL - METHODE II:
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RCPFA_CELL_II IS
    PORT(
        A, B : IN STD_LOGIC;
        FIN, CIN : IN STD_LOGIC;
        FOUT, COUT: OUT STD_LOGIC;
        S : OUT STD_LOGIC
    );
END ENTITY RCPFA_CELL_II;
ARCHITECTURE RCPFA_CELL_II_ARC OF RCPFA_CELL_II IS
    SIGNAL X : STD_LOGIC;
BEGIN
    FOUT <= NOT (A NOR B);
    X <= (A AND B) NOR (NOT CIN);
    S <= X NOR (NOT FIN);
    COUT <= NOT(X NOR NOT(NOT FIN));
END ARCHITECTURE RCPFA_CELL_II_ARC;
-----------------------------------------------------------------------------------
--RFCPA I
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RCPFA_I IS
    PORT(
        A, B : IN STD_LOGIC_VECTOR (15 DOWNTO 0):= (OTHERS=>'0');
        C0: IN STD_LOGIC :='0';
        S : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
END ENTITY RCPFA_I;
ARCHITECTURE RCPFA_I_ARC OF RCPFA_I IS
    SIGNAL F, C : STD_LOGIC_VECTOR (16 DOWNTO 0) := (OTHERS=>'0');
BEGIN
    C(0) <= C0;
    C(16) <= F(16);

     CELL0 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(0), B=>B(0), FIN=>C(0), COUT=>F(0), CIN=>C(1), S=>S(0), FOUT=> F(1));
    CELL1 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(1), B=>B(1), FIN=>F(1), COUT=>C(1), CIN=>C(2), S=>S(1), FOUT=> F(2));
    CELL2 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(2), B=>B(2), FIN=>F(2), COUT=>C(2), CIN=>C(3), S=>S(2), FOUT=> F(3));
    CELL3 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(3), B=>B(3), FIN=>F(3), COUT=>C(3), CIN=>C(4), S=>S(3), FOUT=> F(4));
    CELL4 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(4), B=>B(4), FIN=>F(4), COUT=>C(4), CIN=>C(5), S=>S(4), FOUT=> F(5));
    CELL5 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(5), B=>B(5), FIN=>F(5), COUT=>C(5), CIN=>C(6), S=>S(5), FOUT=> F(6));
    CELL6 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(6), B=>B(6), FIN=>F(6), COUT=>C(6), CIN=>C(7), S=>S(6), FOUT=> F(7));
    CELL7 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(7), B=>B(7), FIN=>F(7), COUT=>C(7), CIN=>C(8), S=>S(7), FOUT=> F(8));
    CELL8 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(8), B=>B(8), FIN=>F(8), COUT=>C(8), CIN=>C(9), S=>S(8), FOUT=> F(9));
    CELL9 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(9), B=>B(9), FIN=>F(9), COUT=>C(9), CIN=>C(10), S=>S(9), FOUT=> F(10));
    CELL19 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(10), B=>B(10), FIN=>F(10), COUT=>C(10), CIN=>C(11), S=>S(10), FOUT=> F(11));
    CELL11 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(11), B=>B(11), FIN=>F(11), COUT=>C(11), CIN=>C(12), S=>S(11), FOUT=> F(12));
    CELL12 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(12), B=>B(12), FIN=>F(12), COUT=>C(12), CIN=>C(13), S=>S(12), FOUT=> F(13));
    CELL13 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(13), B=>B(13), FIN=>F(13), COUT=>C(13), CIN=>C(14), S=>S(13), FOUT=> F(14));
    CELL14 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(14), B=>B(14), FIN=>F(14), COUT=>C(14), CIN=>C(15), S=>S(14), FOUT=> F(15));
    CELL15 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(15), B=>B(15), FIN=>F(15), COUT=>C(15), CIN=>C(16), S=>S(15), FOUT=> F(16));

END ARCHITECTURE RCPFA_I_ARC;

----------------------------------------------------------------------------------
-----------------------------------------------------------------------------------
--RFCPA II
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RCPFA_II IS
    PORT(
        A, B : IN STD_LOGIC_VECTOR (15 DOWNTO 0):= (OTHERS=>'0');
        C0: IN STD_LOGIC :='0';
        S : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
END ENTITY RCPFA_II;
ARCHITECTURE RCPFA_II_ARC OF RCPFA_II IS
    SIGNAL F, C : STD_LOGIC_VECTOR (16 DOWNTO 0) := (OTHERS=>'0');
BEGIN
    C(0) <= C0;
    C(16) <= F(16);

    CELL0 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(0), B=>B(0), FIN=>C(0), COUT=>F(0), CIN=>C(1), S=>S(0), FOUT=> F(1));
    CELL1 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(1), B=>B(1), FIN=>F(1), COUT=>C(1), CIN=>C(2), S=>S(1), FOUT=> F(2));
    CELL2 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(2), B=>B(2), FIN=>F(2), COUT=>C(2), CIN=>C(3), S=>S(2), FOUT=> F(3));
    CELL3 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(3), B=>B(3), FIN=>F(3), COUT=>C(3), CIN=>C(4), S=>S(3), FOUT=> F(4));
    CELL4 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(4), B=>B(4), FIN=>F(4), COUT=>C(4), CIN=>C(5), S=>S(4), FOUT=> F(5));
    CELL5 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(5), B=>B(5), FIN=>F(5), COUT=>C(5), CIN=>C(6), S=>S(5), FOUT=> F(6));
    CELL6 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(6), B=>B(6), FIN=>F(6), COUT=>C(6), CIN=>C(7), S=>S(6), FOUT=> F(7));
    CELL7 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(7), B=>B(7), FIN=>F(7), COUT=>C(7), CIN=>C(8), S=>S(7), FOUT=> F(8));
    CELL8 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(8), B=>B(8), FIN=>F(8), COUT=>C(8), CIN=>C(9), S=>S(8), FOUT=> F(9));
    CELL9 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(9), B=>B(9), FIN=>F(9), COUT=>C(9), CIN=>C(10), S=>S(9), FOUT=> F(10));
    CELL19 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(10), B=>B(10), FIN=>F(10), COUT=>C(10), CIN=>C(11), S=>S(10), FOUT=> F(11));
    CELL11 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(11), B=>B(11), FIN=>F(11), COUT=>C(11), CIN=>C(12), S=>S(11), FOUT=> F(12));
    CELL12 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(12), B=>B(12), FIN=>F(12), COUT=>C(12), CIN=>C(13), S=>S(12), FOUT=> F(13));
    CELL13 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(13), B=>B(13), FIN=>F(13), COUT=>C(13), CIN=>C(14), S=>S(13), FOUT=> F(14));
    CELL14 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(14), B=>B(14), FIN=>F(14), COUT=>C(14), CIN=>C(15), S=>S(14), FOUT=> F(15));
    CELL15 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(15), B=>B(15), FIN=>F(15), COUT=>C(15), CIN=>C(16), S=>S(15), FOUT=> F(16));

END ARCHITECTURE RCPFA_II_ARC;


-----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TB IS
END ENTITY TB;

ARCHITECTURE TEST OF TB IS
    SIGNAL A, B :  STD_LOGIC_VECTOR (15 DOWNTO 0):= (OTHERS=>'0');
    SIGNAL C0:  STD_LOGIC :='0';
    SIGNAL SI, SII :  STD_LOGIC_VECTOR (15 DOWNTO 0);
BEGIN
    CUT_I : ENTITY WORK.RCPFA_I(RCPFA_I_ARC) PORT MAP(A,B,C0,SI);
    CUT_II : ENTITY WORK.RCPFA_II(RCPFA_II_ARC) PORT MAP(A,B,C0,SII);

    A <= X"0001" AFTER 10 NS ,  X"0302" AFTER 30 NS;
    B <= X"0004" AFTER 10 NS ,  X"1009" AFTER 30 NS;

END ARCHITECTURE TEST;



-- FUNCTION G_CALCULATOR ( A_MATRIX ARRAY_TYPE) RETURN ARRAY_TYPE is
-- 	VARIABLE G : STD_LOGIC_VECTOR (7 DOWNTO 0);
-- 	BEGIN
-- 		 FOR I IN O TO 7 LOOP
--             G(I) :=  
-- 	RETURN G;
-- END FUNCTION G_CALCULATOR;




---------------------------------------------------------------------------------------------
-- APROXIMATE HALF ADDER
---------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.std_logic_arith;
ENTITY APPROXIMATE_HALFADDER IS PORT (HALFADDER_INPUT1 : IN STD_LOGIC;
                                        HALFADDER_INPUT2 : IN STD_LOGIC;
                                        HALFADDER_SUM : OUT STD_LOGIC;
                                        HALFADDER_CARRY : OUT STD_LOGIC);
END ENTITY ;

ARCHITECTURE GATE OF APPROXIMATE_HALFADDER IS 
BEGIN 
    HALFADDER_SUM <= HALFADDER_INPUT1 OR HALFADDER_INPUT2;
    HALFADDER_CARRY <= HALFADDER_INPUT1 AND HALFADDER_INPUT2;
END ARCHITECTURE ;

---------------------------------------------------------------------------------------------
-- APROXIMATE FULL ADDER
---------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.std_logic_arith;
ENTITY APPROXIMATE_FULLADDER IS PORT (FULLADDER_INPUT1 : IN STD_LOGIC;
                                        FULLADDER_INPUT2 : IN STD_LOGIC;
                                        FULLADDER_INPUT3 : IN STD_LOGIC;
                                        FULLADDER_SUM : OUT STD_LOGIC;
                                        FULLADDER_CARRY : OUT STD_LOGIC);
END ENTITY ;

ARCHITECTURE GATE OF APPROXIMATE_FULLADDER IS
SIGNAL W : STD_LOGIC;
BEGIN 
    W <= FULLADDER_INPUT1 OR FULLADDER_INPUT2;
    FULLADDER_SUM <= W XOR FULLADDER_INPUT3;
    FULLADDER_CARRY <= W AND FULLADDER_INPUT3;
END ARCHITECTURE; 

---------------------------------------------------------------------------------------------
-- APROXIMATE COMPRESSOR 4 TO 2
---------------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.std_logic_arith;
ENTITY APPROXIMAT_COMPRESSOR4TO2 IS PORT (COMPRESSOR_INPUT1 : IN STD_LOGIC;
                                            COMPRESSOR_INPUT2 : IN STD_LOGIC;
                                            COMPRESSOR_INPUT3 : IN STD_LOGIC;
                                            COMPRESSOR_INPUT4 : IN STD_LOGIC;
                                            COMPRESSOR_SUM : OUT STD_LOGIC;
                                            COMPRESSOR_CARRY : OUT STD_LOGIC);
END ENTITY ;
ARCHITECTURE GATE OF APPROXIMAT_COMPRESSOR4TO2 IS 
SIGNAL W1, W2 : STD_LOGIC;
BEGIN 
    W1 <= COMPRESSOR_INPUT1 AND COMPRESSOR_INPUT2;
    W2 <= COMPRESSOR_INPUT3 AND COMPRESSOR_INPUT4;
    COMPRESSOR_SUM <= (COMPRESSOR_INPUT1 XOR COMPRESSOR_INPUT2) OR (COMPRESSOR_INPUT3 XOR COMPRESSOR_INPUT4) OR (W1 AND W2);
    COMPRESSOR_CARRY <= W1 OR W2;
END ARCHITECTURE;

---------------------------------------------------------------------------------------------
-- Reverse carry propagation full adder
---------------------------------------------------------------------------------------------
--FUNDUMENTAL CELL - METHODE I:
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RCPFA_CELL_I IS
    PORT(
        A, B : IN STD_LOGIC;
        FIN, CIN : IN STD_LOGIC;
        FOUT, COUT: OUT STD_LOGIC;
        S : OUT STD_LOGIC
    );
END ENTITY RCPFA_CELL_I;
ARCHITECTURE RCPFA_CELL_I_ARC OF RCPFA_CELL_I IS
    SIGNAL Y : STD_LOGIC;
BEGIN
    FOUT <= NOT (A NAND B);
    Y <= (A OR B) NAND (NOT CIN);
    S <= Y NAND (NOT FIN);
    COUT <= NOT(Y NAND NOT(NOT FIN));
END ARCHITECTURE RCPFA_CELL_I_ARC;
-----------------------------------------------------------------------------------
--FUNDUMENTAL CELL - METHODE II:
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RCPFA_CELL_II IS
    PORT(
        A, B : IN STD_LOGIC;
        FIN, CIN : IN STD_LOGIC;
        FOUT, COUT: OUT STD_LOGIC;
        S : OUT STD_LOGIC
    );
END ENTITY RCPFA_CELL_II;
ARCHITECTURE RCPFA_CELL_II_ARC OF RCPFA_CELL_II IS
    SIGNAL X : STD_LOGIC;
BEGIN
    FOUT <= NOT (A NOR B);
    X <= (A AND B) NOR (NOT CIN);
    S <= X NOR (NOT FIN);
    COUT <= NOT(X NOR NOT(NOT FIN));
END ARCHITECTURE RCPFA_CELL_II_ARC;
-----------------------------------------------------------------------------------
--RFCPA I
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RCPFA_I IS
    PORT(
        A, B : IN STD_LOGIC_VECTOR (15 DOWNTO 0):= (OTHERS=>'0');
        C0: IN STD_LOGIC :='0';
        S : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
END ENTITY RCPFA_I;
ARCHITECTURE RCPFA_I_ARC OF RCPFA_I IS
    SIGNAL F, C : STD_LOGIC_VECTOR (16 DOWNTO 0) := (OTHERS=>'0');
BEGIN
    C(0) <= C0;
    C(16) <= F(16);

    CELL0 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(0), B=>B(0), FIN=>C(0), COUT=>F(0), CIN=>C(1), S=>S(0), FOUT=> F(1));
    CELL1 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(1), B=>B(1), FIN=>F(1), COUT=>C(1), CIN=>C(2), S=>S(1), FOUT=> F(2));
    CELL2 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(2), B=>B(2), FIN=>F(2), COUT=>C(2), CIN=>C(3), S=>S(2), FOUT=> F(3));
    CELL3 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(3), B=>B(3), FIN=>F(3), COUT=>C(3), CIN=>C(4), S=>S(3), FOUT=> F(4));
    CELL4 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(4), B=>B(4), FIN=>F(4), COUT=>C(4), CIN=>C(5), S=>S(4), FOUT=> F(5));
    CELL5 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(5), B=>B(5), FIN=>F(5), COUT=>C(5), CIN=>C(6), S=>S(5), FOUT=> F(6));
    CELL6 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(6), B=>B(6), FIN=>F(6), COUT=>C(6), CIN=>C(7), S=>S(6), FOUT=> F(7));
    CELL7 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(7), B=>B(7), FIN=>F(7), COUT=>C(7), CIN=>C(8), S=>S(7), FOUT=> F(8));
    CELL8 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(8), B=>B(8), FIN=>F(8), COUT=>C(8), CIN=>C(9), S=>S(8), FOUT=> F(9));
    CELL9 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(9), B=>B(9), FIN=>F(9), COUT=>C(9), CIN=>C(10), S=>S(9), FOUT=> F(10));
    CELL19 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(10), B=>B(10), FIN=>F(10), COUT=>C(10), CIN=>C(11), S=>S(10), FOUT=> F(11));
    CELL11 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(11), B=>B(11), FIN=>F(11), COUT=>C(11), CIN=>C(12), S=>S(11), FOUT=> F(12));
    CELL12 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(12), B=>B(12), FIN=>F(12), COUT=>C(12), CIN=>C(13), S=>S(12), FOUT=> F(13));
    CELL13 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(13), B=>B(13), FIN=>F(13), COUT=>C(13), CIN=>C(14), S=>S(13), FOUT=> F(14));
    CELL14 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(14), B=>B(14), FIN=>F(14), COUT=>C(14), CIN=>C(15), S=>S(14), FOUT=> F(15));
    CELL15 : ENTITY WORK.RCPFA_CELL_I(RCPFA_CELL_I_ARC) PORT MAP(A=>A(15), B=>B(15), FIN=>F(15), COUT=>C(15), CIN=>C(16), S=>S(15), FOUT=> F(16));

END ARCHITECTURE RCPFA_I_ARC;

----------------------------------------------------------------------------------
--RFCPA II
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RCPFA_II IS
    PORT(
        A, B : IN STD_LOGIC_VECTOR (15 DOWNTO 0):= (OTHERS=>'0');
        C0: IN STD_LOGIC :='0';
        S : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
END ENTITY RCPFA_II;
ARCHITECTURE RCPFA_II_ARC OF RCPFA_II IS
    SIGNAL F, C : STD_LOGIC_VECTOR (16 DOWNTO 0) := (OTHERS=>'0');
BEGIN
    C(0) <= C0;
    C(16) <= F(16);

    CELL0 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(0), B=>B(0), FIN=>C(0), COUT=>F(0), CIN=>C(1), S=>S(0), FOUT=> F(1));
    CELL1 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(1), B=>B(1), FIN=>F(1), COUT=>C(1), CIN=>C(2), S=>S(1), FOUT=> F(2));
    CELL2 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(2), B=>B(2), FIN=>F(2), COUT=>C(2), CIN=>C(3), S=>S(2), FOUT=> F(3));
    CELL3 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(3), B=>B(3), FIN=>F(3), COUT=>C(3), CIN=>C(4), S=>S(3), FOUT=> F(4));
    CELL4 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(4), B=>B(4), FIN=>F(4), COUT=>C(4), CIN=>C(5), S=>S(4), FOUT=> F(5));
    CELL5 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(5), B=>B(5), FIN=>F(5), COUT=>C(5), CIN=>C(6), S=>S(5), FOUT=> F(6));
    CELL6 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(6), B=>B(6), FIN=>F(6), COUT=>C(6), CIN=>C(7), S=>S(6), FOUT=> F(7));
    CELL7 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(7), B=>B(7), FIN=>F(7), COUT=>C(7), CIN=>C(8), S=>S(7), FOUT=> F(8));
    CELL8 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(8), B=>B(8), FIN=>F(8), COUT=>C(8), CIN=>C(9), S=>S(8), FOUT=> F(9));
    CELL9 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(9), B=>B(9), FIN=>F(9), COUT=>C(9), CIN=>C(10), S=>S(9), FOUT=> F(10));
    CELL19 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(10), B=>B(10), FIN=>F(10), COUT=>C(10), CIN=>C(11), S=>S(10), FOUT=> F(11));
    CELL11 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(11), B=>B(11), FIN=>F(11), COUT=>C(11), CIN=>C(12), S=>S(11), FOUT=> F(12));
    CELL12 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(12), B=>B(12), FIN=>F(12), COUT=>C(12), CIN=>C(13), S=>S(12), FOUT=> F(13));
    CELL13 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(13), B=>B(13), FIN=>F(13), COUT=>C(13), CIN=>C(14), S=>S(13), FOUT=> F(14));
    CELL14 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(14), B=>B(14), FIN=>F(14), COUT=>C(14), CIN=>C(15), S=>S(14), FOUT=> F(15));
    CELL15 : ENTITY WORK.RCPFA_CELL_II(RCPFA_CELL_II_ARC) PORT MAP(A=>A(15), B=>B(15), FIN=>F(15), COUT=>C(15), CIN=>C(16), S=>S(15), FOUT=> F(16));

END ARCHITECTURE RCPFA_II_ARC;


---------------------------------------------------------------------------------------------
-- complete system_I
---------------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.std_logic_arith;
-- PACKAGE IS
--     TYPE ARRAY_TYPE IS ARRAY OF (NATURAL RANGE <>) STD_LOGIC_VECTOR (7 DOWNTO 0); 
-- END PACKAGE;

ENTITY APPROXIMATE_MULTIPLIER_I IS 
PORT (MULT_INPUT1 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
MULT_INPUT2 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
MULT_OUTPUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END ENTITY ;

ARCHITECTURE GATE OF APPROXIMATE_MULTIPLIER_I IS 

TYPE ARRAY_TYPE IS ARRAY (NATURAL RANGE<>) OF STD_LOGIC_VECTOR(7 DOWNTO 0); 
---CALCULATING "A" USING BOTH INPUT VECTORS:
FUNCTION BITMULTIPLIER (IN1,IN2: STD_LOGIC_VECTOR ) RETURN ARRAY_TYPE IS 
VARIABLE MATRIX : ARRAY_TYPE (7 DOWNTO 0);
BEGIN 
    FOR I IN 0 TO 7 LOOP
        FOR J IN 0 TO 7 LOOP
            MATRIX(I)(J) := IN1(I) AND IN2(J);
        END LOOP;
    END LOOP;
    RETURN MATRIX;
END BITMULTIPLIER;
---------------------------------
-- FUNCTION TO CLACULATE P USING THE A MATRIX
FUNCTION P_CALCULATOR ( A_MATRIX : ARRAY_TYPE) RETURN ARRAY_TYPE is
	VARIABLE P : ARRAY_TYPE (7 DOWNTO 0);
	BEGIN
		 FOR I IN 0 TO 7 LOOP
            FOR J IN 0 TO 7 LOOP
                 P(I)(J) :=  A_MATRIX(I)(J) OR A_MATRIX(J)(I);
            END LOOP;
        END LOOP;
	RETURN P;
END FUNCTION P_CALCULATOR;
---------------------------------
-- FUNCTION TO CLACULATE G USING THE A MATRIX
FUNCTION G_CALCULATOR ( A_MATRIX : ARRAY_TYPE) RETURN ARRAY_TYPE is
	VARIABLE G : ARRAY_TYPE (7 DOWNTO 0);
	BEGIN
		 FOR I IN 0 TO 7 LOOP
            FOR J IN 0 TO 7 LOOP
                 G(I)(J) :=  A_MATRIX(I)(J) AND A_MATRIX(J)(I);
            END LOOP;
        END LOOP;
	RETURN G;
END FUNCTION G_CALCULATOR;

SIGNAL G3, G4, G5, G6, G7, G8, G9, G10, G11 : STD_LOGIC;
SIGNAL S4, S5, S6, S7, S8, S9, S10, S11, S12 : STD_LOGIC;
SIGNAL C4, C5, C6, C7, C8, C9, C10, C11, C12 : STD_LOGIC;
SIGNAL X : STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL Y : STD_LOGIC_VECTOR (15 DOWNTO 0);

SIGNAL G , P, A : ARRAY_TYPE (7 DOWNTO 0);

BEGIN 
-- G3 <= G30 OR G21;
-- G4 <= G40 OR G31;
-- G5 <= G50 OR G41 OR G32;
-- G6 <= G60 OR G51 OR G42;
-- G7 <= G70 OR G61 OR G52 OR G43;
-- G8 <= G71 OR G62 OR G53;
-- G9 <= G72 OR G63 OR G54;
-- G10 <= G73 OR G64;
-- G11 <= G74 OR G65;
A <= BITMULTIPLIER (MULT_INPUT1 , MULT_INPUT2);
P <= P_CALCULATOR (A);
G <= G_CALCULATOR (A);

G3 <= G(3)(0) OR G(2)(1);
G4 <= G(4)(0) OR G(3)(1);
G5 <= G(5)(0) OR G(4)(1) OR G(3)(2);
G6 <= G(6)(0) OR G(5)(1) OR G(4)(2);
G7 <= G(7)(0) OR G(6)(1) OR G(5)(2) OR G(4)(3);
G8 <= G(7)(1) OR G(6)(2) OR G(5)(3);
G9 <= G(7)(2) OR G(6)(3) OR G(5)(4);
G10 <= G(7)(3) OR G(6)(4);
G11 <= G(7)(4) OR G(6)(5);

--FIRST STAGE
HALFADDER1: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (P(4)(0), P(3)(1), S4, C4);
HALFADDER2: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (P(7)(4), P(6)(5), S11, C11);
HALFADDER3: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (A(7)(5), A(5)(7), S12, C12);

FULLADDER1 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(5)(0), P(4)(1), P(3)(2), S5, C5);
FULLADDER2 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(7)(2), P(6)(3), P(5)(4), S9, C9);
FULLADDER3 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(7)(3), P(6)(4), A(5)(5), S10, C10);

COMPRESSOR1 : ENTITY WORK.APPROXIMAT_COMPRESSOR4TO2 PORT MAP (P(6)(0), P(5)(1), P(4)(2), A(3)(3), S6, C6);
COMPRESSOR2 : ENTITY WORK.APPROXIMAT_COMPRESSOR4TO2 PORT MAP (P(7)(0), P(6)(1), P(5)(2), P(4)(3), S7, C7);
COMPRESSOR3 : ENTITY WORK.APPROXIMAT_COMPRESSOR4TO2 PORT MAP (P(7)(1), P(6)(2), P(5)(3), A(4)(4), S8, C8);

--SECOND STAGE
X(0) <= A(0)(0);
Y(0) <= '0';
Y(1) <= '0';

HALFADDER_1: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (A(1)(0), A(0)(1), X(1), Y(2));-- HALFADDER ???

FULLADDER_0 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (A(2)(0), A(0)(2), A(1)(1), X(2), Y(3));
FULLADDER_1 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(3)(0), P(2)(1), G3, X(3), Y(4));
FULLADDER_2 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S4, A(2)(2), G4, X(4), Y(5));
FULLADDER_3 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S5, G5, C4, X(5), Y(6));
FULLADDER_4 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S6, G6, C5, X(6), Y(7));
FULLADDER_5 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S7, G7, C6, X(7), Y(8));
FULLADDER_6 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S8, G8, C7, X(8), Y(9));
FULLADDER_7 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S9, G9, C8, X(9), Y(10));
FULLADDER_8 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S10, G10, C9, X(10), Y(11));
FULLADDER_9 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S11, G11, C10, X(11), Y(12));
FULLADDER_10 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S12, C11, A(6)(6), X(12), Y(13));
FULLADDER_11 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (A(7)(6), A(6)(7), C12, X(13), Y(14));


x(14) <= A(7)(7);

x(15) <= '0';
y(15) <= '0';

--THIRD STAGE 
RCPFA: ENTITY WORK.RCPFA_I PORT MAP (X, Y, '0', MULT_OUTPUT);

END ARCHITECTURE;

---------------------------------------------------------------------------------------------
-- complete system_II
---------------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.std_logic_arith;
-- PACKAGE IS
--     TYPE ARRAY_TYPE IS ARRAY OF (NATURAL RANGE <>) STD_LOGIC_VECTOR (7 DOWNTO 0); 
-- END PACKAGE;

ENTITY APPROXIMATE_MULTIPLIER_II IS 
PORT (MULT_INPUT1 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
MULT_INPUT2 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
MULT_OUTPUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END ENTITY ;

ARCHITECTURE GATE OF APPROXIMATE_MULTIPLIER_II IS 

TYPE ARRAY_TYPE IS ARRAY (NATURAL RANGE<>) OF STD_LOGIC_VECTOR(7 DOWNTO 0); 
---CALCULATING "A" USING BOTH INPUT VECTORS:
FUNCTION BITMULTIPLIER (IN1,IN2: STD_LOGIC_VECTOR ) RETURN ARRAY_TYPE IS 
VARIABLE MATRIX : ARRAY_TYPE (7 DOWNTO 0);
BEGIN 
    FOR I IN 0 TO 7 LOOP
        FOR J IN 0 TO 7 LOOP
            MATRIX(I)(J) := IN1(I) AND IN2(J);
        END LOOP;
    END LOOP;
    RETURN MATRIX;
END BITMULTIPLIER;
---------------------------------
-- FUNCTION TO CLACULATE P USING THE A MATRIX
FUNCTION P_CALCULATOR ( A_MATRIX : ARRAY_TYPE) RETURN ARRAY_TYPE is
	VARIABLE P : ARRAY_TYPE (7 DOWNTO 0);
	BEGIN
		 FOR I IN 0 TO 7 LOOP
            FOR J IN 0 TO 7 LOOP
                 P(I)(J) :=  A_MATRIX(I)(J) OR A_MATRIX(J)(I);
            END LOOP;
        END LOOP;
	RETURN P;
END FUNCTION P_CALCULATOR;
---------------------------------
-- FUNCTION TO CLACULATE G USING THE A MATRIX
FUNCTION G_CALCULATOR ( A_MATRIX : ARRAY_TYPE) RETURN ARRAY_TYPE is
	VARIABLE G : ARRAY_TYPE (7 DOWNTO 0);
	BEGIN
		 FOR I IN 0 TO 7 LOOP
            FOR J IN 0 TO 7 LOOP
                 G(I)(J) :=  A_MATRIX(I)(J) AND A_MATRIX(J)(I);
            END LOOP;
        END LOOP;
	RETURN G;
END FUNCTION G_CALCULATOR;

SIGNAL G3, G4, G5, G6, G7, G8, G9, G10, G11 : STD_LOGIC;
SIGNAL S4, S5, S6, S7, S8, S9, S10, S11, S12 : STD_LOGIC;
SIGNAL C4, C5, C6, C7, C8, C9, C10, C11, C12 : STD_LOGIC;
SIGNAL X : STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL Y : STD_LOGIC_VECTOR (15 DOWNTO 0);

SIGNAL G , P, A : ARRAY_TYPE (7 DOWNTO 0);

BEGIN 
-- G3 <= G30 OR G21;
-- G4 <= G40 OR G31;
-- G5 <= G50 OR G41 OR G32;
-- G6 <= G60 OR G51 OR G42;
-- G7 <= G70 OR G61 OR G52 OR G43;
-- G8 <= G71 OR G62 OR G53;
-- G9 <= G72 OR G63 OR G54;
-- G10 <= G73 OR G64;
-- G11 <= G74 OR G65;
A <= BITMULTIPLIER (MULT_INPUT1 , MULT_INPUT2);
P <= P_CALCULATOR (A);
G <= G_CALCULATOR (A);

G3 <= G(3)(0) OR G(2)(1);
G4 <= G(4)(0) OR G(3)(1);
G5 <= G(5)(0) OR G(4)(1) OR G(3)(2);
G6 <= G(6)(0) OR G(5)(1) OR G(4)(2);
G7 <= G(7)(0) OR G(6)(1) OR G(5)(2) OR G(4)(3);
G8 <= G(7)(1) OR G(6)(2) OR G(5)(3);
G9 <= G(7)(2) OR G(6)(3) OR G(5)(4);
G10 <= G(7)(3) OR G(6)(4);
G11 <= G(7)(4) OR G(6)(5);

--FIRST STAGE
HALFADDER1: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (P(4)(0), P(3)(1), S4, C4);
HALFADDER2: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (P(7)(4), P(6)(5), S11, C11);
HALFADDER3: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (A(7)(5), A(5)(7), S12, C12);

FULLADDER1 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(5)(0), P(4)(1), P(3)(2), S5, C5);
FULLADDER2 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(7)(2), P(6)(3), P(5)(4), S9, C9);
FULLADDER3 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(7)(3), P(6)(4), A(5)(5), S10, C10);

COMPRESSOR1 : ENTITY WORK.APPROXIMAT_COMPRESSOR4TO2 PORT MAP (P(6)(0), P(5)(1), P(4)(2), A(3)(3), S6, C6);
COMPRESSOR2 : ENTITY WORK.APPROXIMAT_COMPRESSOR4TO2 PORT MAP (P(7)(0), P(6)(1), P(5)(2), P(4)(3), S7, C7);
COMPRESSOR3 : ENTITY WORK.APPROXIMAT_COMPRESSOR4TO2 PORT MAP (P(7)(1), P(6)(2), P(5)(3), A(4)(4), S8, C8);

--SECOND STAGE
X(0) <= A(0)(0);
Y(0) <= '0';
Y(1) <= '0';

HALFADDER_1: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (A(1)(0), A(0)(1), X(1), Y(2));-- HALFADDER ???

FULLADDER_0 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (A(2)(0), A(0)(2), A(1)(1), X(2), Y(3));
FULLADDER_1 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(3)(0), P(2)(1), G3, X(3), Y(4));
FULLADDER_2 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S4, A(2)(2), G4, X(4), Y(5));
FULLADDER_3 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S5, G5, C4, X(5), Y(6));
FULLADDER_4 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S6, G6, C5, X(6), Y(7));
FULLADDER_5 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S7, G7, C6, X(7), Y(8));
FULLADDER_6 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S8, G8, C7, X(8), Y(9));
FULLADDER_7 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S9, G9, C8, X(9), Y(10));
FULLADDER_8 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S10, G10, C9, X(10), Y(11));
FULLADDER_9 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S11, G11, C10, X(11), Y(12));
FULLADDER_10 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S12, C11, A(6)(6), X(12), Y(13));
FULLADDER_11 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (A(7)(6), A(6)(7), C12, X(13), Y(14));


x(14) <= A(7)(7);

x(15) <= '0';
y(15) <= '0';

--THIRD STAGE 
RCPFA: ENTITY WORK.RCPFA_II PORT MAP (X, Y, '0', MULT_OUTPUT);

END ARCHITECTURE;





---------------------------------------------------------------------------------------------
-- complete system CLA
---------------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.std_logic_arith;
-- PACKAGE IS
--     TYPE ARRAY_TYPE IS ARRAY OF (NATURAL RANGE <>) STD_LOGIC_VECTOR (7 DOWNTO 0); 
-- END PACKAGE;

ENTITY APPROXIMATE_MULTIPLIER_CPA IS 
PORT (MULT_INPUT1 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
MULT_INPUT2 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
MULT_OUTPUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END ENTITY ;

ARCHITECTURE GATE OF APPROXIMATE_MULTIPLIER_CPA IS 

TYPE ARRAY_TYPE IS ARRAY (NATURAL RANGE<>) OF STD_LOGIC_VECTOR(7 DOWNTO 0); 
---CALCULATING "A" USING BOTH INPUT VECTORS:
FUNCTION BITMULTIPLIER (IN1,IN2: STD_LOGIC_VECTOR ) RETURN ARRAY_TYPE IS 
VARIABLE MATRIX : ARRAY_TYPE (7 DOWNTO 0);
BEGIN 
    FOR I IN 0 TO 7 LOOP
        FOR J IN 0 TO 7 LOOP
            MATRIX(I)(J) := IN1(I) AND IN2(J);
        END LOOP;
    END LOOP;
    RETURN MATRIX;
END BITMULTIPLIER;
---------------------------------
-- FUNCTION TO CLACULATE P USING THE A MATRIX
FUNCTION P_CALCULATOR ( A_MATRIX : ARRAY_TYPE) RETURN ARRAY_TYPE is
	VARIABLE P : ARRAY_TYPE (7 DOWNTO 0);
	BEGIN
		 FOR I IN 0 TO 7 LOOP
            FOR J IN 0 TO 7 LOOP
                 P(I)(J) :=  A_MATRIX(I)(J) OR A_MATRIX(J)(I);
            END LOOP;
        END LOOP;
	RETURN P;
END FUNCTION P_CALCULATOR;
---------------------------------
-- FUNCTION TO CLACULATE G USING THE A MATRIX
FUNCTION G_CALCULATOR ( A_MATRIX : ARRAY_TYPE) RETURN ARRAY_TYPE is
	VARIABLE G : ARRAY_TYPE (7 DOWNTO 0);
	BEGIN
		 FOR I IN 0 TO 7 LOOP
            FOR J IN 0 TO 7 LOOP
                 G(I)(J) :=  A_MATRIX(I)(J) AND A_MATRIX(J)(I);
            END LOOP;
        END LOOP;
	RETURN G;
END FUNCTION G_CALCULATOR;

SIGNAL G3, G4, G5, G6, G7, G8, G9, G10, G11 : STD_LOGIC;
SIGNAL S4, S5, S6, S7, S8, S9, S10, S11, S12 : STD_LOGIC;
SIGNAL C4, C5, C6, C7, C8, C9, C10, C11, C12 : STD_LOGIC;
SIGNAL X : STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL Y : STD_LOGIC_VECTOR (15 DOWNTO 0);

SIGNAL G , P, A : ARRAY_TYPE (7 DOWNTO 0);

BEGIN 
-- G3 <= G30 OR G21;
-- G4 <= G40 OR G31;
-- G5 <= G50 OR G41 OR G32;
-- G6 <= G60 OR G51 OR G42;
-- G7 <= G70 OR G61 OR G52 OR G43;
-- G8 <= G71 OR G62 OR G53;
-- G9 <= G72 OR G63 OR G54;
-- G10 <= G73 OR G64;
-- G11 <= G74 OR G65;
A <= BITMULTIPLIER (MULT_INPUT1 , MULT_INPUT2);
P <= P_CALCULATOR (A);
G <= G_CALCULATOR (A);

G3 <= G(3)(0) OR G(2)(1);
G4 <= G(4)(0) OR G(3)(1);
G5 <= G(5)(0) OR G(4)(1) OR G(3)(2);
G6 <= G(6)(0) OR G(5)(1) OR G(4)(2);
G7 <= G(7)(0) OR G(6)(1) OR G(5)(2) OR G(4)(3);
G8 <= G(7)(1) OR G(6)(2) OR G(5)(3);
G9 <= G(7)(2) OR G(6)(3) OR G(5)(4);
G10 <= G(7)(3) OR G(6)(4);
G11 <= G(7)(4) OR G(6)(5);

--FIRST STAGE
HALFADDER1: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (P(4)(0), P(3)(1), S4, C4);
HALFADDER2: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (P(7)(4), P(6)(5), S11, C11);
HALFADDER3: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (A(7)(5), A(5)(7), S12, C12);

FULLADDER1 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(5)(0), P(4)(1), P(3)(2), S5, C5);
FULLADDER2 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(7)(2), P(6)(3), P(5)(4), S9, C9);
FULLADDER3 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(7)(3), P(6)(4), A(5)(5), S10, C10);

COMPRESSOR1 : ENTITY WORK.APPROXIMAT_COMPRESSOR4TO2 PORT MAP (P(6)(0), P(5)(1), P(4)(2), A(3)(3), S6, C6);
COMPRESSOR2 : ENTITY WORK.APPROXIMAT_COMPRESSOR4TO2 PORT MAP (P(7)(0), P(6)(1), P(5)(2), P(4)(3), S7, C7);
COMPRESSOR3 : ENTITY WORK.APPROXIMAT_COMPRESSOR4TO2 PORT MAP (P(7)(1), P(6)(2), P(5)(3), A(4)(4), S8, C8);

--SECOND STAGE
X(0) <= A(0)(0);
Y(0) <= '0';
Y(1) <= '0';

HALFADDER_1: ENTITY WORK.APPROXIMATE_HALFADDER PORT MAP (A(1)(0), A(0)(1), X(1), Y(2));-- HALFADDER ???

FULLADDER_0 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (A(2)(0), A(0)(2), A(1)(1), X(2), Y(3));
FULLADDER_1 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (P(3)(0), P(2)(1), G3, X(3), Y(4));
FULLADDER_2 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S4, A(2)(2), G4, X(4), Y(5));
FULLADDER_3 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S5, G5, C4, X(5), Y(6));
FULLADDER_4 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S6, G6, C5, X(6), Y(7));
FULLADDER_5 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S7, G7, C6, X(7), Y(8));
FULLADDER_6 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S8, G8, C7, X(8), Y(9));
FULLADDER_7 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S9, G9, C8, X(9), Y(10));
FULLADDER_8 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S10, G10, C9, X(10), Y(11));
FULLADDER_9 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S11, G11, C10, X(11), Y(12));
FULLADDER_10 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (S12, C11, A(6)(6), X(12), Y(13));
FULLADDER_11 : ENTITY WORK.APPROXIMATE_FULLADDER PORT MAP (A(7)(6), A(6)(7), C12, X(13), Y(14));


x(14) <= A(7)(7);

x(15) <= '0';
y(15) <= '0';

--THIRD STAGE 
CPA: ENTITY WORK.CPA_n PORT MAP (X, Y, '0', MULT_OUTPUT);

END ARCHITECTURE;




